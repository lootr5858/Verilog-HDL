module  c_tb();

reg		clk;
reg		rst;
reg		en;

wire [7:0] val;
wire		  reached;

